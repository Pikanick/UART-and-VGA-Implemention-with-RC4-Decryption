library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity lab3 is
    port(
        CLOCK_50            : in  std_logic;
        KEY                 : in  std_logic_vector(3 downto 0);
        SW                  : in  std_logic_vector(17 downto 0);
        VGA_R, VGA_G, VGA_B : out std_logic_vector(9 downto 0);  -- The outs go to VGA controller
        VGA_HS              : out std_logic;
        VGA_VS              : out std_logic;
        VGA_BLANK           : out std_logic;
        VGA_SYNC            : out std_logic;
        VGA_CLK             : out std_logic
    );
end lab3;

architecture rtl of lab3 is

 --Component from the Verilog file: vga_adapter.v

    component vga_adapter
        generic(RESOLUTION : string);
        port (
            resetn                                          : in  std_logic;
            clock                                           : in  std_logic;
            colour                                          : in  std_logic_vector(2 downto 0);
            x                                               : in  std_logic_vector(7 downto 0);
            y                                               : in  std_logic_vector(6 downto 0);
            plot                                            : in  std_logic;
            VGA_R, VGA_G, VGA_B                             : out std_logic_vector(9 downto 0);
            VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_CLK    : out std_logic
        );
    end component;

    component line_drawer is
        port(
            clk_i       : in std_logic;
            rst_i       : in std_logic;
    
            colour_o    : out std_logic_vector(2 downto 0);
            x_o         : out std_logic_vector(7 downto 0);
            y_o         : out std_logic_vector(6 downto 0);
            plot_o      : out std_logic
        );
    end component;

    signal colour       : std_logic_vector(2 downto 0);
    signal plot         : std_logic;
    signal x            : std_logic_vector(7 downto 0);
    signal y            : std_logic_vector(6 downto 0);

    signal rst_active_1 : std_logic;

begin

  -- includes the vga adapter, which should be in your project

    rst_active_1 <= not KEY(3);

    vga_u0 : vga_adapter
        generic map(RESOLUTION => "160x120")
        port map(
            resetn    => KEY(3),
            clock     => CLOCK_50,
            colour    => colour,
            x         => x,
            y         => y,
            plot      => plot,
            VGA_R     => VGA_R,
            VGA_G     => VGA_G,
            VGA_B     => VGA_B,
            VGA_HS    => VGA_HS,
            VGA_VS    => VGA_VS,
            VGA_BLANK => VGA_BLANK,
            VGA_SYNC  => VGA_SYNC,
            VGA_CLK   => VGA_CLK
        );

    line_drawer0 : line_drawer
        port map(
            clk_i       => CLOCK_50,
            rst_i       => rst_active_1,
            colour_o    => colour,
            x_o         => x,
            y_o         => y,
            plot_o      => plot
        );

end architecture;

